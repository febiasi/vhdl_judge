-- Teste


Lets see...
